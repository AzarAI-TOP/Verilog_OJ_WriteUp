module P1 (
    output one
);
  // Write your code here
  assign one = 1'b1;
endmodule
