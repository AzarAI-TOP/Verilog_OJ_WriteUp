module P3 (
    input  in,
    output out
);
  // Write your code here
  assign out = in;
endmodule
