module P6 (
    input  a,
    input  b,
    output out
);
  // 请用户在下方编辑代码
  assign out = a & b;

  //用户编辑到此为止
endmodule
