module P2 (
    output out
);
  // Write your code here
  assign out = 1'b0;
endmodule
