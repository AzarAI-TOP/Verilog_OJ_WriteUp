module P4 (
    input a,
    input b,
    input c,

    output w,
    output x,
    output y,
    output z
);
  // write your code below
  assign w = a;
  assign x = b;
  assign y = b;
  assign z = c;

endmodule
