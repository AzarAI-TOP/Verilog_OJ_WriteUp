module P5 (
    input  in,
    output out
);
  // write your code below
  assign out = ~in;
endmodule
